//Interface
interface dut_if1;

//Input signals
logic a_in;
logic b_in;
logic c_in;

//Output_signals
logic sum_out;
logic carry_out;

//Control Signals
logic clock;
logic reset;

endinterface
