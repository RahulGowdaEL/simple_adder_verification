//SEQR

class adder_seqr extends uvm_sequencer;
`uvm_component_utils(adder_seqr)

function new(string name = adder_seqr, uvm_component parent);
   super.new(name,parent);
endfunction
endclass
